module mux_8x1_tb;
  reg [2:0] s1;
  reg [7:0] i1;
  reg [7:0] y1;
  
  mux_8x1 m8 (.i(i1), .s(s1), .y(y1));
  
  initial begin
    $dumpfile("dump.vcd");
    $dumpvars();
    $monitor("time=%0t, i1=%d, s1=%b, y1=%d", $time, i1, s1, y1);
    
    
    #5 {s1[2], s1[1], s1[0]} = 3'b000; i1 = 8'b00000001;
    #5 {s1[2], s1[1], s1[0]} = 3'b001; i1 = 8'b00000010;
    #5 {s1[2], s1[1], s1[0]} = 3'b010; i1 = 8'b00000100;
    #5 {s1[2], s1[1], s1[0]} = 3'b011; i1 = 8'b00001000;
    #5 {s1[2], s1[1], s1[0]} = 3'b100; i1 = 8'b00010000;
    #5 {s1[2], s1[1], s1[0]} = 3'b101; i1 = 8'b00100000;
    #5 {s1[2], s1[1], s1[0]} = 3'b110; i1 = 8'b01000000;
    #5 {s1[2], s1[1], s1[0]} = 3'b111; i1 = 8'b10000000;
    
    #10 $finish;
  end
endmodule
