// Code your testbench here
// or browse Examples

module all_logic_gates_tb;
  
  reg a,b;
  wire not_gate,
       and_gate,
       or_gate,
       nand_gate,
       nor_gate,
       xor_gate,
       xnor_gate;
  
  all_logic_gates dut(a,b,not_gate,and_gate,or_gate,nand_gate,nor_gate,xor_gate,xnor_gate);
  
  initial
    begin
      
      $dumpfile("dump.vcd");
      $dumpvars(0,all_logic_gates_tb);
      
            $monitor("time=%0t,a=%b,b=%b,not_gate=%0d,and_gate=%0d,or_gate=%0d,nand_gate=%0d,nor_gate=%0d,xor_gate=%0d,xnor_gate= %0d",$time,a,b,not_gate,and_gate,or_gate,nand_gate,nor_gate,xor_gate,xnor_gate);

      // for all 4 states
      #1 a = 1'b0; b = 1'b0;
      #1 a = 1'b0; b = 1'b1;
      #1 a = 1'b0; b = 1'bx;
      #1 a = 1'b0; b = 1'bz;
      
      // for all 4 states

      #1 a = 1'b1; b = 1'b0;
      #1 a = 1'b1; b = 1'b1;
      #1 a = 1'b1; b = 1'bx;
      #1 a = 1'b1; b = 1'bz;
      
      // for all 4 states

      #1 a = 1'bx; b = 1'b0;
      #1 a = 1'bx; b = 1'b1;
      #1 a = 1'bx; b = 1'bx;
      #1 a = 1'bx; b = 1'bz;
      
      // for all 4 states
      
      #1 a = 1'bz; b = 1'b0;
      #1 a = 1'bz; b = 1'b1;
      #1 a = 1'bz; b = 1'bx;
      #1 a = 1'bz; b = 1'bz;
      
      #30;
      $finish;
    end
endmodule
      
  